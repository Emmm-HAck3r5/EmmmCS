`define YAMM_IDLE 0
`define YAMM_1BYTE 1
`define YAMM_2BYTE 2
`define YAMM_3BYTE 3
`define YAMM_4BYTE 4
`define YAMM_FINISHED 5

`define YAMM_VGA_MEM_OPR 6
`define YAMM_VGA_REG_OPR 7
`define YAMM_LED_OPR 8
`define YAMM_MEM_OPR 9

`define YAMM_VGA_MEM_OPR_FIN 10
`define YAMM_VGA_MEM_REG_FIN 11
`define YAMM_LED_OPR_FIN 12
`define YAMM_1BYTE_FIN 13
`define YAMM_2BYTE_FIN 14
`define YAMM_3BYTE_FIN 15
`define YAMM_4BYTE_FIN 16

`define YAMM_MODE_R32 0
`define YAMM_MODE_W8 1
`define YAMM_MODE_W16 2
`define YAMM_MODE_W32 3

`define YAMM_MEM 0
`define YAMM_VGA_MEM 1
`define YAMM_LED_MEM 2

//hard coded
`define YAMM_MEM_BEGIN 32'h0
`define YAMM_MEM_END 32'h80000
`define YAMM_VGA_MEM_BEGIN 32'h80004
`define YAMM_VGA_MEM_END 32'h812C4
`define YAMM_VGA_REG_BEGIN 32'h812C4
`define YAMM_VGA_REG_END 32'h812C6
`define YAMM_LED_MEM_BEGIN 32'h80000
`define YAMM_LED_MEM_END 32'h80002

//hard coded
`define YAMM_LED_ADDR1 32'h80000
`define YAMM_LED_ADDR2 32'h80001
`define YAMM_VGA_CURSOR_X 32'h812C4
`define YAMM_VGA_CURSOR_Y 32'h812C5
module cpu_bus(
	input 						clk,
	input						reset_n,
	input	[31:0]				address,
	input	[31:0]				wdata,
	input	[1:0]				WLEN,
	input						EN_N,
	output reg					READY,
	output reg [31:0]			rdata,
	// debugging
	output 			global_wen,
	output			cache_en,
	output			cache_wen,
	output reg [15:0] selected_rdata,
	output reg  [31:0] addr_offset,
	output reg [2:0]	bus_state,
	output wire [15:0] cache_rdata,
	output reg [15:0] wdata16,
	output wire [31:0] vgac_addr,
	/////////////// LED ///////////////
	output 			[9:0]		LEDR,
	/////////////// VGA ///////////////
	output		          		VGA_BLANK_N,
	output		    [7:0]		VGA_B,
	output		          		VGA_CLK,
	output		    [7:0]		VGA_G,
	output		          		VGA_HS,
	output		    [7:0]		VGA_R,
	output		          		VGA_SYNC_N,
	output		          		VGA_VS
);

`define ADDR_SIZE		32
`define WORD_SIZE		16
`define BYTE_SIZE		8

`define	CACHE_MAXSIZE	32'h80000
`define	LED_MAXSIZE		32'h4
`define VGA_MEMORY_SIZE	32'h12C0
`define VGA_CREGS_SIZE  32'h10

`define	CACHE_START		32'h0
`define	LED_START		(`CACHE_START + `CACHE_MAXSIZE)
`define	VGA_START		(`LED_START + `LED_MAXSIZE)
`define VGA_CTRL_START	(`VGA_START + `VGA_MEMORY_SIZE)
`define	KB_START		(`VGA_CTRL_START + `VGA_CREGS_SIZE)

// ENABLE
// wire cache_en;
wire led_en;
wire vga_en;
wire vgac_en;
assign cache_en = (address >= `CACHE_START) && (address < `LED_START);
assign led_en = (address >= `LED_START) && (address < `VGA_START);
assign vga_en =  (address >= `VGA_START) && (address < `VGA_CTRL_START);
assign vgac_en =  (address >= `VGA_CTRL_START) && (address < `KB_START);

// base ADDRESS
wire [`ADDR_SIZE - 1:0] cache_addr;
wire [`ADDR_SIZE - 1:0] led_addr;
wire [`ADDR_SIZE - 1:0] vga_addr;
// wire [`ADDR_SIZE - 1:0] vgac_addr;
wire [`ADDR_SIZE - 1:0] vga_dp_raddr;
// reg  [`ADDR_SIZE - 1:0] addr_offset;

assign cache_addr = address - `CACHE_START + addr_offset;
assign led_addr = address - `LED_START + addr_offset;
assign vga_addr = address - `VGA_START + addr_offset;
assign vgac_addr = address - `VGA_CTRL_START + addr_offset;

// select output radata
// wire [`WORD_SIZE - 1:0] cache_rdata;
wire [`WORD_SIZE - 1:0] led_rdata;
wire [`WORD_SIZE - 1:0] vga_rdata;
wire [`WORD_SIZE - 1:0] vgac_rdata;
wire [`WORD_SIZE - 1:0] vga_dp_rdata;
// reg [`WORD_SIZE - 1:0] selected_rdata;

always @ (negedge clk)
	if (cache_en) selected_rdata <= cache_rdata;
	else if (led_en) selected_rdata <= led_rdata;
	else if (vga_en) selected_rdata <= vga_rdata;
	else if (vgac_en) selected_rdata <= vgac_rdata;
	else selected_rdata <= selected_rdata;

// write-in data
// wire global_wen;
// wire cache_wen;
wire led_wen;
wire vga_wen;
wire vgac_wen;
// reg [`WORD_SIZE - 1:0] wdata16;
reg writing = 0;

assign global_wen = writing;
assign cache_wen = cache_en && global_wen;
assign led_wen = led_en && global_wen;
assign vga_wen = vga_en && global_wen;
assign vgac_wen = vgac_en && global_wen;

// ADDRESS MAPPING FSM
`define BUS_ST_IDLE			0
`define	BUS_ST_RD32_R1		1
`define	BUS_ST_RD32_R2		2
`define	BUS_ST_WR8_R		3
`define	BUS_ST_WR8_W		4
`define	BUS_ST_WR16_W		5
`define	BUS_ST_WR32_W1		6
`define	BUS_ST_WR32_W2		7

`define WLEN_RD32	2'b00
`define WLEN_WR8	2'b01
`define WLEN_WR16	2'b10
`define WLEN_WR32	2'b11

// reg [2:0] bus_state = `BUS_ST_IDLE;

initial begin
	bus_state = `BUS_ST_IDLE;
end

// address offset
always @ (posedge clk) begin
	case (bus_state)
	  `BUS_ST_IDLE:
	  	if (!EN_N && WLEN == `WLEN_RD32)
		  addr_offset <= 32'd2;
		else addr_offset <= 32'd0;
	  `BUS_ST_WR32_W1: addr_offset <= 32'd2;
	  default: addr_offset <= 32'd0;
	endcase
end

// select read data
always @ (posedge clk) begin
	case (bus_state)
	  `BUS_ST_RD32_R1: rdata[`WORD_SIZE-1:0] <= selected_rdata;
	  `BUS_ST_RD32_R2: rdata[2*`WORD_SIZE-1:`WORD_SIZE] <= selected_rdata;
	  default: rdata <= rdata;
	endcase
end

// writing
always @ (posedge clk)
	case (bus_state)
		`BUS_ST_WR8_W, `BUS_ST_WR16_W, `BUS_ST_WR32_W2: writing <= 0;
		`BUS_ST_WR8_R: writing <= 1;
		`BUS_ST_IDLE:
			if (!EN_N)
				case (WLEN)
					`WLEN_RD32, `WLEN_WR8: writing <= 0;
					`WLEN_WR16, `WLEN_WR32: writing <= 1;
				endcase
			else writing <= 0;
		default: writing <= writing;
	endcase

// write-in data
always @ (posedge clk) begin
	case(bus_state)
		`BUS_ST_WR8_R:
			if (address[0]) wdata16 <= {wdata[7:0], selected_rdata[7:0]};
			else wdata16 <= {selected_rdata[`WORD_SIZE-1:8], wdata[7:0]};
		`BUS_ST_WR32_W1:  wdata16 <= wdata[2*`WORD_SIZE-1:`WORD_SIZE];
		default: wdata16 <= wdata[`WORD_SIZE-1:0];
	endcase
end

// state transformation
always @ (posedge clk) begin
	case (bus_state)
		`BUS_ST_IDLE : begin
			READY <= 1;
			if (EN_N) bus_state <= `BUS_ST_IDLE;
			else begin
				READY <= 0;
				case (WLEN)
					`WLEN_RD32: bus_state <= `BUS_ST_RD32_R1;
					`WLEN_WR8: bus_state <= `BUS_ST_WR8_R;
					`WLEN_WR16: bus_state <= `BUS_ST_WR16_W;
					`WLEN_WR32: bus_state <= `BUS_ST_WR32_W1;
				  	default: bus_state <= `BUS_ST_IDLE;
				endcase
			end
		end
		`BUS_ST_RD32_R1:bus_state <= `BUS_ST_RD32_R2;
		`BUS_ST_RD32_R2:bus_state <= `BUS_ST_IDLE;
		`BUS_ST_WR8_R:bus_state <= `BUS_ST_WR8_W;
		`BUS_ST_WR8_W:bus_state <= `BUS_ST_IDLE;
		`BUS_ST_WR16_W:bus_state <= `BUS_ST_IDLE;
		`BUS_ST_WR32_W1:bus_state <= `BUS_ST_WR32_W2;
		`BUS_ST_WR32_W2:bus_state <= `BUS_ST_IDLE;
	  default: bus_state <= `BUS_ST_IDLE;
	endcase
end

// MEMORYS
reg [`WORD_SIZE - 1 : 0] led_memory [(`LED_MAXSIZE / 2) - 1 : 0];
reg [`VGA_CREGS_SIZE * `BYTE_SIZE - 1 : 0 ] vga_ctrl = 0;

cache c(
	.address(cache_addr[18:1]),
	.clock(clk),
	.data(wdata16),
	.wren(cache_wen),
	.q(cache_rdata)
	);

vga_memory2port vm2p(
	.clock(clk),
	// display ctrl only read
	.address_a(vga_dp_raddr[11:0]),
	// data_a is not used
	.wren_a(0),
	.q_a(vga_dp_rdata),
	// vga memory write/read
	.address_b(vga_addr[12:1]),
	.data_b(wdata16),
	.wren_b(vga_wen),
	.q_b(vga_rdata)
);

assign led_rdata = led_memory[0];

always @ (posedge clk) begin
	if (led_wen && address[1:0] < 2'b10) begin
		led_memory[led_addr[1]] <= wdata16;
	end
end

reg [`WORD_SIZE - 1 : 0] vgac_save;
assign vgac_rdata = vgac_save;
initial vga_ctrl = 0;
always @ (posedge clk) begin
	if (~vgac_addr[4])
		vgac_save <= vga_ctrl[{vgac_addr[3:1], 4'hf} -: `WORD_SIZE];
	else vgac_save <= 16'h0;
	if (vgac_wen && ~vgac_addr[4]) begin
		// MAGIC OPERATORS '+:' / '-:'
		vga_ctrl[{vgac_addr[3:1], 4'hf} -: `WORD_SIZE] <= wdata16;
	end
end

// DEVICE OUTPUT
assign LEDR = led_memory[0][9:0];

wire [7:0] x_addr;
wire [4:0] y_addr;

assign vga_dp_raddr = ({7'b0,y_addr} << 6) + ({7'b0,y_addr} << 4) + x_addr;

display_ctrl dp(
    .clk(clk),
    .reset_n(reset_n),
    .in_data(vga_dp_rdata),
    .ctrl_reg(vga_ctrl),
    .x_addr(x_addr),
    .y_addr(y_addr),
    .vga_rst(~reset_n),
    .vga_vs(VGA_VS),
    .vga_hs(VGA_HS),
    .vga_syncn(VGA_SYNC_N),
    .vga_blankn(VGA_BLANK_N),
    .vga_clk(VGA_CLK),
    .vga_r(VGA_R),
    .vga_g(VGA_G),
    .vga_b(VGA_B)
    );

endmodule
