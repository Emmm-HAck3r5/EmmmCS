/*
  Copyright 2018 EmmmHackers

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

        http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
  --------------------------
  File: cpu_gregs.v
  Project: EmmmCS
  File Created: 2018-11-20 23:19:54
  Author: Chen Haodong (easyai@outlook.com)
  --------------------------
  Last Modified: 2018-11-21 16:30:19
  Modified By: Chen Haodong (easyai@outlook.com)
 */

`include "cpu_define.v"

module cpu_gregs(
    input clk,
    input rd_wen,

    input [`CPU_GREGIDX_WIDTH-1:0] rs1_idx,
    input [`CPU_GREGIDX_WIDTH-1:0] rs2_idx,
    input [`CPU_GREGIDX_WIDTH-1:0] rd_idx,

    output reg [`CPU_XLEN-1:0] rs1_dat,
    output reg [`CPU_XLEN-1:0] rs2_dat,
    input [`CPU_XLEN-1:0] rd_dat
    );
    reg [`CPU_XLEN-1:0] rx [`CPU_GREG_COUNT-1:0];

    always @(posedge clk)
    begin
        rx[0] = `CPU_XLEN'b0;
        rs1_dat = rx[rs1_idx];
        rs2_dat = rx[rs2_idx];
        if(rd_wen && rd_idx!=`CPU_GREGIDX_WIDTH'b0)
        begin
            rx[rd_idx] = rd_dat;
        end
    end
endmodule